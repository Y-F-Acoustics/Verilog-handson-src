module mydivider_2(CLK_i, CLK_o);
    /*
        mydivider.v
        clock divider (dividing ratio: 1/2)

        // port definition
        Input
        -----
            CLK_i : Input clock

        Output
        ------
            CLK_o : Output divided clock
    */

    /* Port definition */
    // Input
    input wire CLK_i;

    // Output
    output wire CLK_o;

    /* Internal Register */
    // Write register definition if you need

    /* RTL */
    // Write your code here

endmodule