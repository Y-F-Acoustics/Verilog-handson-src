module combfilter(CLK_i, data_in, data_out);
    /*
		  combfilter.v
      combfilter

      // Port definition
      Input
      -----
        CLK_i : input clock
        data_in : 4 bit input data

      Output
      ------
        CLK_o : output clock
        data_out : output data
    */

    /* Port definition */
    // Input
    /* Write input port definition here */

    // Output
    /* Write input port definition here */

    /* Register definition */
    /* Write internal register definition here if you need */

    /* RTL */
    /* Write your code here */
    
endmodule