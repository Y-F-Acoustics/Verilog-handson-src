module mycounter_4bit(CLK, out);
    /*
		mycounter_4bit.v
        4 bit counter with clock

        // Port definition
        Input
        -----
            CLK: counter clock

        Output
        ------
            out: 4 bit unsigned integer increments with positive edge  of clock
    */

    /* Port definition */
    // Input
    /* write input definition here */

    // Output
    /* write output definition here */

    /* Internal register */
    /* write internal register here if you need */

    /* RTL */
    always @ (/*Write Sensitivity List Here*/) begin
        /* Write your code here */
    end


endmodule