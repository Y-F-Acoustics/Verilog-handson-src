module FullAdder(A, B, C, out, cy);
/*
  FullAdder.v
    1 bit Full Adder.

    // Port Definition
    Input
    -----
        A, B, C: 1 bit input number

    Output
    ------
        out: 1 bit Result
        cy : Carry bit
*/

/* Port Definition */
// Inputs
/* Write your code here to meet port definition */

// Outputs
output wire out;
output wire cy; 

/* Internal Signal Definition (If you need) */
/* Write code here if you need */

/* RTL */
/* Write your code here to meet specification */

endmodule