`timescale 1 us/ 1 ns
module test_mycounter();
    /*
        test_mycounter.v
        test bench for mycounter_4bit

        // Signal definition
        in_CLK: input for CLK
        out_out: output for out
    */

    /* Signal definition */
    /* Input signal definition here */

    /* Instantiation */
    /* Write Instantiation here */

    /* Generate clock */
    always begin
        #10 /* Write your test code here */
    end
endmodule