module HalfAdder(A, B, out, cy);
/*
  HalfAdder.v
    1 bit Half Adder.

    // Port Definition
    Input
    -----
        A, B: 1 bit input number

    Output
    ------
        out: 1 bit Result
        cy : Carry bit
*/

/* Port definition */
// Inputs
input wire A, B;

// Outputs
output wire out;
output wire cy;


/* Internal Signal definition (If you need) */
// Write internal signal here if you need.


/* RTL */
// Write circuit description here.

endmodule